entity b is
  port(e1,e2 : in bit;
       f: out bit);
end b;

architecture arch1 of b is
begin
end arch1;

architecture arch2 of b is
begin
end arch2;
